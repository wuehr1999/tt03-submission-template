`timescale 1ns/10ps

module test_top (
    input wire [7:0] io_in,
    output wire [7:0] io_out
);

endmodule
